module reg_file #(
    parameter WIDTH = 32
) (
    input logic ad1,
    input logic ad2,
    input logic ad3,
    input logic we3,
    input logic wd3,
    input logic clk,
    output logic rd1,
    output logic rd2,
    output logic a0
);
endmodule
