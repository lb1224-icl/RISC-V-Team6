module control_unit #(
    
) (
    input logic                    imm_src,
    input logic  [11:0]            imm,
    output logic [WIDTH-1:0]  imm_op
);

endmodule 
