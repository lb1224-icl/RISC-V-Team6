module reg_file #(
    parameter
    D_WIDTH = 8,
    A_WIDTH = 8
) (
    input logic ad1,
    input logic ad2,
    input logic ad3,
    input logic we3,
    input logic wd3,
    input logic clk,
    output logic rd1,
    output logic rd2,
    output logic a0
);
endmodule
